module not_gate_behav(a, y);
  input a;
  output y;
  assign y = ~a;
endmodule