module demux1to4_behav (
  input data_in,      
  input [1:0] sel,    
  output reg [3:0] out
);

  always @(*) begin
    
    out = 4'b0000; 
    
    case (sel)
      2'b00: out[0] = data_in; // Se sel=00, out[0] recebe o dado
      2'b01: out[1] = data_in; // Se sel=01, out[1] recebe o dado
      2'b10: out[2] = data_in; // Se sel=10, out[2] recebe o dado
      2'b11: out[3] = data_in; // Se sel=11, out[3] recebe o dado
    endcase
  end

endmodule